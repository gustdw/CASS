module testbench;
initial begin
    $display("Your SystemVerilog simulator works!");
    $finish;
end
endmodule




